module Elevator(clk32Hz,)

